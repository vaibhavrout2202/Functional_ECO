module patch (g2, g1, t_0);
	input g2, g1;
	output t_0;
	or (t_0, g1, g2);


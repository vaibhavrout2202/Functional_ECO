module patch(t_0, g2, g1);
	input g2, g1;
	output t_0;
	or (t_0, g1, g2);
endmodule
